//-----------------------------------------------------------------------------------------------------------------
//ReadMe: 
// Top module for testing purposes.
// This file (TOP.v) is intended to test the first step of integration between
// UART communication and PSRAM external memory. The test protocol is the following:

// STEP ONE - Initialization: RGB LEDs will start off. By pressing Button B,
// the PSRAM initialization will start. When LEDs turn white, it means PSRAM was
// successfully initialized and it is on its idle state.

// STEP TWO - After initialization, MSGA will be written to PSRAM.
// NOTE: From this step forward, Button B needs to be pressed in order to move
// to next step

// STEP THREE -   MSGA will be read from PSRAM. Upon pressing Button B, stored
// message will be sent through UART. Also, the script will move to next step

// STEP FOUR - Message was also stored to a local reg. Press Button A to sweep
// through the saved data.

// STEP FIVE ONWARDS - Same as STEP TWO, THREE AND FOUR, for MSGB.

// NOTES: 
// Upon error, RED LED will be displayed. 
// During debugging, blue light will turn on
// During process, green led will turn on
//-----------------------------------------------------------------------------------------------------------------

//Include sub-modules (SIMULATION ONLY)
//`include "PSRAM.v" //Simulation modules
//`include "gowin_rpll/grPLL_27_to_84.v" //rPLL Gowin native module


//-----------------------------------------------------------------------------------------------------------------
// TOP MODULE
module TOP (

//Tang Nano 1k
input sys_clk,                //Internal 27 MHz oscillator
input buttonA,                //Tang Nano Button A
input buttonB,                //Tang Nano Button B

//UART
input uart_rx,                 //RX UART wire pin 18

//PSRAM mem chip
inout [3:0] mem_sio,     // sio[0] pin 40, sio[1] pin 39, sio[2] pin 38, sio[3] pin 41
output mem_ce,                // pin 42
output mem_clk_enabled,             // pin 6
output uart_tx,                // TX UART wire pin 17

//DEBUGGING
//Debug RGB LED
output reg [2:0] led_rgb     //RGB LEDs

//Debug external LEDs
//output reg [3:0] led
);

//-----------------------------------------------------------------------------------------------------------------
//Variables

//Wire

//UART-PSRAM interface
reg [22:0] address;       //Address of message to be written/read
//wire [15:0] message;

wire [15:0] write;
reg send_uart;


wire quad_start_uart;         //Start reading OR writing proccess via UART
wire [1:0] read_write_uart;   //Read or write switch via UART
wire [22:0] address_uart;     //Address of interest (write or read) via UART
wire [15:0] data_in_uart;     //Data to be written via UART


//Button A synchronisation and debouncing
wire buttonA_debounced;
//Button B synchronisation and debouncing
wire buttonB_debounced;

//PSRAM interface
wire [15:0] data_out;      //Data read -> Output reg from PSRAM

//Reg
//PSRAM interface
reg [15:0] data_in;         //Data to be written (16 bits)
reg [15:0] read;            //Auxiliary Data read -> reg to be changed at procedural script
reg error;                  //Error flag
reg quad_start;            // Flag to start QPI communication
reg d_com_start;
reg com_start;
// Debugging
reg [3:0] process; //Keep track of write and reading test processes
reg [3:0] counter; //Counter to control debugging LEDs when pressing buttonA
reg [1:0] read_write;
reg pause;

//Directly control write and read process, through MCU (Gowin)
reg [1:0] read_write_mcu;
reg quad_start_mcu;
reg [22:0] address_mcu;
reg [15:0]debug;
reg [15:0] data_in_mcu;

//-----------------------------------------------------------------------------------------------------------------

//SUBMODULES

//84Mhz generated by Gowin's PLL
gowin_rpll_27_to_84 clk2(
    .clkout(clk_PSRAM), //84 MHz
    .clkin(sys_clk) //27MHz
);

//Debouncing processes to avoid noise from button pressing
//sync_debouncer debuttonA(
//    .clk(clk_PSRAM),
//    .button(buttonA),
//    .button_once(buttonA_debounced)
//);

sync_debouncer debuttonB(
    .clk(clk_PSRAM),
    .button(buttonB),
    .button_once(buttonB_debounced)
);

//PSRAM initialization
psram initialize(
    //input
    .mem_clk(clk_PSRAM),
    .startbu(buttonB_debounced),
    .address(address),
    .read_write(read_write),
    .data_in(data_in),
    .quad_start(quad_start),

    //output
    .mem_clk_enabled(mem_clk_enabled),
    .qpi_on(qpi_on),
    .endcommand(endcommand),
    .mem_ce(mem_ce),
    .data_out(data_out),

    //inout
    .mem_sio(mem_sio)
    //.message(message)
);

//UART1 channel communication
uart #(.DELAY_FRAMES(234), .BUFFER_LENGTH(BUFFER_LENGTH)) UART1 (
    //input
    .sys_clk(sys_clk),
    .uart_rx(uart_rx),
    .send_msg(read),
    .send_uart(send_uart),
    
    //output
    .read_write(read_write_uart),
    .quad_start(quad_start_uart),
    .data_in(data_in_uart),
    //.message(message),
    .address(address_uart),
    .uart_tx(uart_tx)
);

//-----------------------------------------------------------------------------------------------------------------

//LOCAL PARAMETERS

//Testbench read & write
localparam [3:0] WRITE_MCU_INIT = 0;
localparam [3:0] READ_MCU_INIT = 1;
localparam [3:0] CHECK_STARTUP = 2;
localparam [3:0] IDLE = 3;
localparam [3:0] WRITE_MCU = 4;
localparam [3:0] READ_MCU = 5;

//CHANGING PARAMETERS
//localparam [15:0] ADDRESSA = 16'h01;
//localparam [15:0] ADDRESSB = 16'h01;
//localparam [15:0] MSGA = 16'h0121;
//localparam [15:0] MSGB = 16'h0123;

//Number of bytes stored in buffer
localparam BUFFER_LENGTH = 6;

//-----------------------------------------------------------------------------------------------------------------

//SCRIPT
initial begin
    process <= WRITE_MCU_INIT;
    error <= 0;
    counter <= 0;
    pause <= 0;
    read <= 0;
    send_uart <= 0;
    com_start <= 0;
    d_com_start <= 0;
    debug <= 0;

    //MCU read-write variables
    read_write_mcu <= 0;
    read_write_mcu <= 0;
    address_mcu <= 0;
    data_in_mcu <= 0;
end



always @(quad_start_mcu || quad_start_uart) begin
    if (process == IDLE) begin
        read_write = read_write_uart;
        address = address_uart;
        data_in = data_in_uart;
        quad_start = quad_start_uart;
    end else begin
        read_write = read_write_mcu;
        address = address_mcu;
        data_in = data_in_mcu;
        quad_start = quad_start_mcu;
    end
end

always @(posedge clk_PSRAM) begin

    d_com_start <= com_start;

    //Detect a rising edge of mcu requisition. Only valid on MCU controlling of WRITE/READs
    quad_start_mcu <= (com_start && ~d_com_start);
    
    //Testing PSRAM communication
    if (qpi_on) begin  //if on IDLE state

      //White LED to begin process
      led_rgb[2:0] <= 3'b000;

      //LED RGBs
      if(error) led_rgb[2:0] <= 3'b011;           //Red LED
      else if (process == WRITE_MCU_INIT || process == READ_MCU_INIT) led_rgb[2:0] <= 3'b010;    //Blue LED = debugging state
      else if (process == IDLE) led_rgb[2:0] <= 3'b101;
      else led_rgb[2:0] <= 3'b000;

      send_uart <= 0;   //Reset send_uart to only be triggered once. Subject to changes
        
        case(pause)

          0: begin
            case (process)

              WRITE_MCU_INIT: begin

                address_mcu <= 24'hABCD;
                data_in_mcu <= 16'h1234;
                read_write_mcu <= 1;
                com_start <= 1;

                if(endcommand) begin
                  debug <= 1;
                  com_start <= 0;
                  process <= READ_MCU_INIT;
                end
              end

              READ_MCU_INIT: begin

                read_write_mcu <= 2;
                com_start <= 1;

                if(endcommand) begin
                  read <= data_out;
                  process <= CHECK_STARTUP;
                  read_write_mcu <= 0;
                  com_start <= 0;
                end
              end

              CHECK_STARTUP: begin
                if(read == data_in_mcu) begin
                  debug <= read;
                  led_rgb <= 3'b101;
                  error <= 0;
                  process <= IDLE;
                end
                else begin
                  error <= 1;
                end
             end
              
              //Writing operation
              IDLE: begin
                if(endcommand && read_write == 2) begin   //Se uma leitura tiver sido requisitada e endcommand = 1..
                    process <= WRITE_MCU;
                    read <= data_out;
                    send_uart <= 1;           // Flag para enviar mensagem na UART
                end
                else if(endcommand && read_write == 1) begin   //Se uma escrita tiver sido requisitada e endcommand = 1..
                    process <= READ_MCU;
                    //send_uart <= 1;           // Flag para enviar mensagem na UART
                end
              end

            WRITE_MCU: begin

                address_mcu <= 24'hABCD;
                data_in_mcu <= 16'h1234;
                read_write_mcu <= 1;

                com_start <= 1;

                if(endcommand) begin
                  process <= IDLE;
                  read_write_mcu <= 0;
                  com_start <= 0;
                end
              end

              READ_MCU: begin
                address_mcu <= 24'h1234;
                read_write_mcu <= 2;
                com_start <= 1;

                if(endcommand) begin
                  process <= IDLE;
                  read <= data_out;
                  read_write_mcu <= 0;
                  com_start <= 0;
                end
              end
            endcase
          end
    
          1: begin //Awaits for button pressed
            if(buttonB_debounced) begin
                pause <= 0;
                //process <= process + 1;
            end
          end

        endcase
      end
end

endmodule

