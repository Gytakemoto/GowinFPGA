//ReadMe: Top module for simulation purposes. To simulate in Icarus Verilog, inside Tang-Nano-1k/src type in cmd:
//iverilog -o Testbench.vvp Testbench.v
//vvp Testbench.vvp
//gtkwave.exe .\Testbench.vcd
//Refer to TOP.V for testing purposes
//----------------------------------------------------------------------------------------------------------------------

//Include sub-modules
`include "PSRAM_simu.v" //Simulation modules
`include "gowin_rpll/grPLL_27_to_84.v" //rPLL Gowin native module

`timescale 1us/1fs
module Testbench ();

//Variables

//Clock varibles
wire sys_clk;             //Internal clock 27MHz
wire clk_PSRAM;         //PSRAM clock 84 MHz
reg enable;            //Clock enable

//Initialization variables
reg startbutton;            //Start when button is pressed
wire [3:0] step;            //Step of initialization
wire [3:0] mem_sio;         //SIO[3:0] ports
wire [15:0] timer;          //Time counter
wire mem_ce;                //PSRAM chip enable
wire [7:0] command;
reg [23:0] address;        //Address of message to be written/read
reg write_sw;
reg read_sw;
reg [15:0] data_in; 
wire [15:0] data_out;
reg [3:0] estepe; //APAGAR depois
reg error;
reg go;
reg [15:0] read;
wire [5:0] counter;


//Clock generation

//27MHz (simulates internal clock)
clk_gen clk1(
    .enable(enable),
    .clk(sys_clk)
);

//84Mhz generated by Gowin's PLL
Gowin_rPLL_27_to_84MHz clk2(
    .clkout(clk_PSRAM), //84 MHz
    .clkin(sys_clk) //27MHz
);

//PSRAM initialization
psram_simu initialize(
    //input
    .mem_clk(clk_PSRAM),
    .startbu(startbutton),
    .address(address),
    .read_sw(read_sw),
    .write_sw(write_sw),
    .data_in(data_in),

    //output
    .counter(counter),
    .endcommand(endcommand),
    .mem_ce(mem_ce),
    .step(step),
    .command(command),
    .data_out(data_out),

    //inout
    .mem_sio(mem_sio)
);

parameter real PSRAM_FREQ = 84;
parameter real clk_pd = 1/(PSRAM_FREQ * 1e6) * 1e9;

//Testbench read & write
localparam [3:0] WRITEA = 0;
localparam [3:0] WRITEB = 1;
localparam [3:0] READA = 2;
localparam [3:0] READB = 3;
localparam [3:0] NEXT = 4;

initial begin
    estepe <= 0;
    error <= 0;
end

always @(posedge clk_PSRAM) begin
    if (go)
      begin
        case (estepe)
          WRITEA: begin   
            address <= 8'h12;
            data_in <= 16'h1234;
            write_sw <= 1;
            if(endcommand) begin
               estepe <= WRITEB;
               write_sw <= 0;
            end
          end
          WRITEB: begin   
            address <= 8'h2;
            data_in <= 16'h5678;
            write_sw <= 1;
            if(endcommand) begin
              estepe <= READA;
              write_sw <= 0;
            end
          end
          READA: begin
            address <= 8'h12;
            read_sw <= 1;
            if(endcommand) begin 
              estepe <= READB;
              read_sw <= 0;
            end
          end
          READB: begin
            read <= data_out;
            if ( data_out != 16'h1234 ) begin   
              error <= 1;            
            end
            address <= 8'h2;
            read_sw <= 1;
            if(endcommand) begin 
              estepe <= NEXT;
              read_sw <= 0;
            end
          end
          NEXT: begin
            read <= data_out;
            if ( data_out != 16'h3456 ) begin 
              error <= 1;
            end
            //if(endcommand) estepe <= WRITEA;
          end        
        endcase     
      end
end

//Proccess simulation
initial begin
    //$display ("PSRAM desired FREQ: %0.3f ns", clk_pd);
    $dumpfile("Testbench.vcd");
    $dumpvars(1, Testbench);

    write_sw = 0;
    read_sw = 0;
    go = 0;
    error = 0;

    #50 enable = 1;
    #100 startbutton = 1;

    //Write proccess
    #500 go = 1;


    #500 startbutton = 0;
    enable = 0;

    $finish; 
end

endmodule
