
/* ------------------------------- TOP MODULE ------------------------------- */
module TOP (

//Tang Nano 1k
input sys_clk,                	// Internal 27 MHz oscillator

//UART
input uart_rx,                 	// RX UART wire [pin 18]

//PSRAM mem chip
inout [3:0] mem_sio,     		// Communication busbar for PSRAM communication - [sio[0] pin 40, sio[1] pin 39, sio[2] pin 38, sio[3] pin 41]
output mem_ce,                	// PSRAM chip enable - [pin 42]
output mem_clk_enabled,         // PSRAM clock pin - [pin 6]
output uart_tx,                	// TX UART wire [pin 17]

//DEBUGGING
//Debug RGB LED
output reg [2:0] led_rgb,     	// RGB LEDs

//Debug external LEDs
output [3:0] led				// Debugs external LEDs
);

/* -------------------------------- Variables ------------------------------- */

/* ----------------------------- PSRAM interface ---------------------------- */

// Inputs (from PSRAM.v module)
wire clk_PSRAM;				   // 84MHz rPLL generated clock. Used in PSRAM interface
wire endcommand;			   // Input flag - indicates whether PSRAM writing or reading finished
wire qpi_on;				   // Input flag - indicates whether QPI communication is on

// Outputs (to PSRAM.v module) - Determined by "MCU" or UART
reg [22:0] address;       	   // Address of message to be written/read
reg [15:0] data_in;            // Data to be written (16 bits)
reg [15:0] read;               // Auxiliary Data read -> reg receives data_out in a procedural script
wire [15:0] data_out;      	   // Data read -> Output reg from PSRAM
reg [1:0] read_write;		   // Define read or write proccess
	//read_write
	//0	0 : Do nothing
	//0	1 : Write data from PSRAM
    //1	0 : Read data to PSRAM
    //1	1 : Do nothing


/* ----------------------------- UART interface ----------------------------- */

// Inputs (from UART.v module)
	// Request read or write through UART
wire quad_start_uart;         // Start reading OR writing proccess via UART
wire [1:0] read_write_uart;   // Read or write switch via UART
wire [22:0] address_uart;     // Address of interest (write or read) via UART
wire [15:0] data_in_uart;     // Data to be written via UART

// Outputs (to UART.v module)
reg send_uart;				  // Flag - inform UART to send data through Tx

/* -------------------------- Internal variables -------------------------- */

reg error;                  // Error flag
reg [3:0] process; 			// State-machine of top.v states

// Request read or write through MCU
reg com_start;				// Detect rising edge to start quad_start
reg d_com_start;			
reg quad_start;            	// Output flag - Start reading OR writing proccess via MCU
	// quad_start = com_start && !d_com_start;

// Directly control write and read process, through MCU (Gowin)
reg quad_start_mcu;
reg [1:0] read_write_mcu;
reg [22:0] address_mcu;
reg [15:0] data_in_mcu;

/* ------------------------------- Submodules ------------------------------- */

/* --------------------- 84Mhz generated by Gowin's PLL --------------------- */
gowin_rpll_27_to_84 clk2(
	.clkout(clk_PSRAM), 	// 84 MHz
	.clkin(sys_clk) 		// 27MHz
);

/* ---------------------------------- PSRAM --------------------------------- */
psram initialize(
	//input
	.mem_clk(clk_PSRAM),
	.address(address),
	.read_write(read_write),
	.data_in(data_in),
	.quad_start(quad_start),

	//output
	.mem_clk_enabled(mem_clk_enabled),
	.qpi_on(qpi_on),
	.endcommand(endcommand),
	.mem_ce(mem_ce),
	.data_out(data_out),

	//inout
	.mem_sio(mem_sio)
);

/* ----------------------- UART1 channel communication ---------------------- */
uart #(.DELAY_FRAMES(729), .BUFFER_LENGTH(BUFFER_LENGTH)) UART1 (
	//input
	.clk_PSRAM(clk_PSRAM),
	.uart_rx(uart_rx),
	.send_msg(read),
	.send_uart(send_uart),
	
	//output
	.led(led),
	.read_write(read_write_uart),
	.quad_start(quad_start_uart),
	.data_in(data_in_uart),
	.address(address_uart),
	.uart_tx(uart_tx)
);

/* ---------------------------- Local parameters ---------------------------- */

//Testbench read & write
localparam [3:0] WRITE_MCU_INIT = 0;
localparam [3:0] READ_MCU_INIT = 1;
localparam [3:0] CHECK_STARTUP = 2;
localparam [3:0] IDLE = 3;

//Buffer's bytes length
localparam BUFFER_LENGTH = 6;

/* --------------------------- Procedural routine --------------------------- */

initial begin
	process <= WRITE_MCU_INIT;
	error <= 0;
	read <= 0;
	send_uart <= 0;
	com_start <= 0;
	d_com_start <= 0;

	//MCU read-write variables
	read_write_mcu <= 0;
	address_mcu <= 22'hzzzz;
	data_in_mcu <= 0;
	quad_start_mcu <= 0;
    led_rgb <= 3'b111;
end

always @(posedge clk_PSRAM) begin

	//* Constantly update regulators in order to avoid inferred latches
	quad_start <= 0;
	read_write <= read_write;
	address <= address;
	data_in <= data_in;
	read <= read;
	send_uart <= 0;

	// Detect a rising edge of mcu requisition. Only valid on MCU controlling of WRITE/READs
	quad_start_mcu <= (com_start && ~d_com_start);
	d_com_start <= com_start;
	com_start <= 0;

    // Routine to detect source of requisition: UART or MCU
	if(quad_start_mcu || quad_start_uart) begin
		//! UART only works while at IDLE state
		if (process == IDLE) begin
			read_write <= read_write_uart;
			address <= address_uart;
			data_in <= data_in_uart;
			quad_start <= quad_start_uart;
		end else begin
			read_write <= read_write_mcu;
			address <= address_mcu;
			data_in <= data_in_mcu;
			quad_start <= quad_start_mcu;
		end
	end

	//* Only when QPI is ready
	if (qpi_on) begin
		case (process)
		    // Writing operation to test PSRAM before starting
			WRITE_MCU_INIT: begin
				address_mcu <= 24'hABCD;
				data_in_mcu <= 16'h1234;
				read_write_mcu <= 1;
				com_start <= 1;
				if(endcommand) begin
					com_start <= 0;
					process <= READ_MCU_INIT;
				end
			end
			READ_MCU_INIT: begin
				address_mcu <= 24'hABCD;
				read_write_mcu <= 2;
				com_start <= 1;
				if(endcommand) begin
					read <= data_out;
					read_write_mcu <= 0;
					com_start <= 0;
					process <= CHECK_STARTUP;
				end
			end
			CHECK_STARTUP: begin
				//* If writing and reading processess were OK
				if(read == data_in_mcu) begin
					led_rgb <= 3'b101;
					error <= 0;
					process <= IDLE;
				end
				// If not...
				else begin
                    led_rgb[2:0] <= 3'b011;
					error <= 1;
				end
			end
			// Writing operation
			IDLE: begin
				if (endcommand) begin
					
					// Read operation
					if (read_write == 2) begin
						read <= data_out;
                        send_uart <= 1;  // Flag to send message via UART
					end
					// Write operation
					else if (read_write == 1) begin
						read <= data_in;
                        send_uart <= 1;  // Flag to send message via UART
					end
                    // Change RGB LED colors
                    if(led_rgb[2:0] == 3'b111) begin
						led_rgb[2:0] <= 3'b000;
                    end 
                    else begin
						led_rgb[2:0] <= {led_rgb[2:0] + 3'd1};  // +1 per LED update
                    end
				end
				process <= IDLE;
			end
		endcase
	end
end
endmodule

