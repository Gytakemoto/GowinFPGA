//ReadMe: Top module for testing purposes.
//Refer to Testbench.v for simulation purposes
//PSRAM communication WITH the need to state beginning and ending of communication. Choosen architecture due to future work (fingers crossed)
//-----------------------------------------------------------------------------------------------------------------

//Include sub-modules
//`include "PSRAM.v" //Simulation modules
//`include "gowin_rpll/grPLL_27_to_84.v" //rPLL Gowin native module

module TOP (

//IO pins
//INPUT
input sys_clk, //Internal 27 MHz oscillator
input buttonA, //Tang Nano Button A
input buttonB, //Tang Nano Button B

//PSRAM mem chip
inout [3:0] mem_sio,    // sio[0] pin 40, sio[1] pin 39, sio[2] pin 38, sio[3] pin 41
output mem_ce,               // pin 42
output mem_clk_en,            // pin 6

//OUTPUT
//Debug RGB LED
output reg [2:0] led_rgb,             //RGB LEDs

//Debug external LEDs
output reg [3:0] led
);

//Variables
//Write/read variables
wire [15:0] message;        //inout variable responsible to send and receive commands to be written and readen, respectively

//Reg

//PSRAM communication
reg [23:0] address;         //Address of message to be written/read
reg [15:0] msg_reg = 0;     //Reg variable of message used in procedural assignment
reg com_start;             //Flag indicates whether start QPI or not
reg d_com_start;
wire quad_start;
reg [1:0] read_write;               //Read enable switch
//  R   W   RW
//  0   0   0   :   Idle state
//  0   1   1   :   Writintg
//  1   0   2   :   Reading
//  1   1   3   :   Undefined


//DEBUGGING
reg [15:0] read;            //Auxiliary Data read -> reg to be changed at procedural script -> debug LEDs
reg error;                  //Error flag
reg [3:0] counter;          //Counter to control debugging LEDs when pressing buttonA
reg pause;                  //Pause flag in order to debug. Proccess MUST work without pauses
reg [3:0] debug_main;

//TOP operation
reg [3:0] proccess;         //Keep track of write and reading test proccesses
reg [15:0] data_in;
wire [15:0] data_out;


//When sending a message, assumes data in msg_reg (msg_uart)
//assign message = (read_write == 1) ? msg_reg:16'hz;

assign quad_start = (com_start & ~d_com_start);

//Button A synchronisation and debouncing
wire buttonA_debounced;

//Button B synchronisation and debouncing
wire buttonB_debounced;

//84Mhz generated by Gowin's PLL
gowin_rpll_27_to_84 clk2(
    .clkout(clk_PSRAM), //84 MHz
    .clkin(sys_clk) //27MHz
);


//Debouncing proccesses to avoid noise from button pressing
sync_debouncer debuttonA(
    .clk(clk_PSRAM),
    .button(buttonA),
    .button_once(buttonA_debounced)
);

sync_debouncer debuttonB(
    .clk(clk_PSRAM),
    .button(buttonB),
    .button_once(buttonB_debounced)
);

//PSRAM initialization
psram initialize(
    //input
    .mem_clk(clk_PSRAM),
    .startbu(buttonB),
    .address(address),
    .read_write(read_write),
    .quad_start(quad_start),
    .data_in(data_in),

    //output
    .mem_clk_en(mem_clk_en),
    .qpi_on(qpi_on),
    .endcommand(endcommand),
    .mem_ce(mem_ce),
    .data_out(data_out),

    //inout
    .mem_sio(mem_sio),
    .message(message)
);

//Testbench read & write
localparam [3:0] WRITEA = 0;
localparam [3:0] WRITEB = 1;
localparam [3:0] READA = 2;
localparam [3:0] READB = 3;
localparam [3:0] WAITA = 4;
localparam [3:0] WAITB = 5;

//CHANGING PARAMETERS
//localparam [22:0] ADDRESSA = 23'h7FFFFF;
localparam [22:0] ADDRESSA = 23'h7FFFFE;
localparam [15:0] ADDRESSB = 16'hABCD;
localparam [15:0] MSGA = 16'h1234;
localparam [15:0] MSGB = 16'h4464;


initial begin
    proccess <= 0;
    error <= 0;
    counter <= 0;
    pause <= 0;
    read_write <= 0;
    com_start <= 0;
    d_com_start <= 0;
    debug_main<= 0;
    read <= 16'hffff;
    address <= 22'h0000;
end

always @(posedge clk_PSRAM) begin

    d_com_start <= com_start;

   //Activates only when error is present while pressing buttonA
   if((error || proccess == WAITA || proccess == WAITB) && buttonA_debounced) begin

        counter <= counter + 1'd1;

        //For each button pressed, change debug LEDs
        case(counter) 
            0: led[3:0] <= read[15:12];
            1: led[3:0] <= read[11:8];
            2: led[3:0] <= read[7:4];
            3: led[3:0] <= read[3:0];
            4: begin
                led[3:0] <= 4'b1111;
                counter <= 0;

            end
            default: begin
                counter <= 0;
            end
        endcase
    end

    //White LED to begin debugging
    led_rgb[2:0] <= 3'b000;

    //Testing PSRAM communication
    if (qpi_on) begin  //if on IDLE state

      //LED RGBs
      if(error) led_rgb[2:0] <= 3'b011;           //Red LED
      else if ((proccess == WAITA || proccess == WAITB)) led_rgb[2:0] <= 3'b110;    //Blue LED = waiting state
      else if ((proccess == WRITEA || proccess == WRITEB)) led_rgb[2:0] <= 3'b010;    //Purple LED = writing state
      else if ((proccess == READA || proccess == READB)) led_rgb[2:0] <= 3'b001;    //Yellow LED = reading state
      else led_rgb[2:0] <= 3'b111;    //LEDs off = Idle, awaiting button
      
      //Keep regs updated
      read <= read;
      com_start <= com_start;
      ////proccess <= proccess;
      address <= address;

        case(pause)

          0: begin
            case (proccess)

              //Writing operation
              WRITEA: begin 
                address <= ADDRESSA;
                data_in <= MSGA;
                //msg_reg <= MSGA;

                //Start writing communication
                read_write <= 1;
                com_start <= 1;
                //pause <= 0;

                if(endcommand) begin
                    proccess <= READA;
                    //Stop communication
                    com_start <= 0;
                    //pause <= 1;
                end
              end

              //Reading operation
              READA: begin
                address <= ADDRESSA;
                //Start reading communication
                read_write <= 2;
                com_start <= 1;

                if(endcommand) begin
                  read <= data_out;
                  debug_main <= 1'd1;
                  //Stop communication
                  com_start <= 0;
                  proccess <= WAITA;
                  //pause <= 1;
                  //read <= message;
                end
              end

              //Awaits for instructions
               WAITA: begin   
                 if ( read == MSGA ) begin   
                    error <= 0; 
                  end
                  else error <= 1;
                  //proccess <= WRITEB;
               end

              //Writing operation
              WRITEB: begin   
                address <= ADDRESSB;
                //msg_reg <= MSGB;
                data_in <= MSGB;
                read_write <= 1;
                com_start <= 1;
                if(endcommand) begin
                    proccess <= READB;
                    com_start <= 0;
                    //pause <= 1;
                end
              end

              //Reading proccess
              READB: begin
                address <= ADDRESSB;
                read_write <= 2;
                com_start <= 1;
                if(endcommand) begin
                  read <= data_out; 
                  com_start <= 0;
                  proccess <= WAITB;
                  //pause <= 1;
                  //read <= message;
                end
              end

              //Awaits for instructions
              WAITB: begin   
                 if ( read == MSGB && !error) begin   
                    error <= 0;
                    led_rgb[2:0] <= 3'b101;     //Comms' succeeded
                  end
                  else error <= 1;
               end
            endcase    
          end

          1: begin //Awaits for button pressed
            if(buttonB_debounced) pause <= 0;
          end

        endcase
      end
end

endmodule

