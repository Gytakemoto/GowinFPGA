//Include sub-modules
`include "PSRAM_simu.v" //Simulation modules
`include "gowin_rpll/grPLL_27_to_84.v" //rPLL Gowin native module

`timescale 1us/1fs
module Testbench ();

//Variables

//Clock varibles
wire clock;             //Internal clock 27MHz
wire clk_PSRAM;         //PSRAM clock 84 MHz
reg enable;            //Clock enable

//Initialization variables
reg startbutton;            //Start when button is pressed
wire [3:0] step;            //Step of initialization
wire [3:0] mem_sio;  //SIO[3:0] ports
wire [15:0] timer;          //Time counter
wire mem_ce;                //PSRAM chip enable
wire [7:0] command;

//Clock generation

//27MHz (simulates internal clock)
clk_gen clk1(
    .enable(enable),
    .clk(clock)
);

//84Mhz generated by Gowin's PLL
Gowin_rPLL_27_to_84MHz clk2(
    .clkout(clk_PSRAM), //84 MHz
    .clkin(clock) //27MHz
);

//PSRAM initialization
psram initialize(
    .sys_clk(clock),
    .mem_clk(clk_PSRAM),
    .startbu(startbutton),
    .mem_sio(mem_sio),
    .mem_ce(mem_ce),
    .step(step),
    .timer(timer),
    .command(command)
);

parameter real PSRAM_FREQ = 84;
parameter real clk_pd = 1/(PSRAM_FREQ * 1e6) * 1e9;


//Proccess simulation
initial begin
    //$display ("PSRAM desired FREQ: %0.3f ns", clk_pd);
    $dumpfile("Testbench.vcd");
    $dumpvars(1, Testbench);
    #200 enable = 1;
    #300 startbutton = 1;

    #500 startbutton = 0;
    enable = 0;

    $finish; 
end

endmodule
