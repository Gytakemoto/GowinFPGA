module onoff (
    input btn_i,
    output led //011 -> Green color
);

assign led = btn_i;

endmodule