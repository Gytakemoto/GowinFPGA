//-----------------------------------------------------------------------------------------------------------------
//ReadMe: 
// Top module for testing purposes.
// This file (TOP.v) is intended to test the first step of integration between
// UART communication and PSRAM external memory. The test protocol is the following:

// STEP ONE - Initialization: RGB LEDs will start off. By pressing Button B,
// the PSRAM initialization will start. When LEDs turn white, it means PSRAM was
// successfully initialized and it is on its idle state.

// STEP TWO - After initialization, MSGA will be written to PSRAM.
// NOTE: From this step forward, Button B needs to be pressed in order to move
// to next step

// STEP THREE -   MSGA will be read from PSRAM. Upon pressing Button B, stored
// message will be sent through UART. Also, the script will move to next step

// STEP FOUR - Message was also stored to a local reg. Press Button A to sweep
// through the saved data.

// STEP FIVE ONWARDS - Same as STEP TWO, THREE AND FOUR, for MSGB.

// NOTES: 
// Upon error, RED LED will be displayed. 
// During debugging, blue light will turn on
// During proccess, green led will turn on
//-----------------------------------------------------------------------------------------------------------------

//Include sub-modules (SIMULATION ONLY)
//`include "PSRAM.v" //Simulation modules
//`include "gowin_rpll/grPLL_27_to_84.v" //rPLL Gowin native module


//-----------------------------------------------------------------------------------------------------------------
// TOP MODULE
module TOP (

//Tang Nano 1k
input sys_clk,                //Internal 27 MHz oscillator
input buttonA,                //Tang Nano Button A
input buttonB,                //Tang Nano Button B

//UART
input uart_rx,                 //RX UART wire pin 18

//PSRAM mem chip
inout [3:0] mem_sio,     // sio[0] pin 40, sio[1] pin 39, sio[2] pin 38, sio[3] pin 41
output mem_ce,                // pin 42
output clk_PSRAM,             // pin 6
output uart_tx,                // TX UART wire pin 17

//DEBUGGING
//Debug RGB LED
output reg [2:0] led_rgb,     //RGB LEDs

//Debug external LEDs
output reg [3:0] led
);

//-----------------------------------------------------------------------------------------------------------------
//Variables

//Wire

//UART-PSRAM interface
wire [23:0] address;
wire [15:0] message;
wire read_psram;
wire read_uart;
wire write_uart;
reg [15:0] write;


//Button A synchronisation and debouncing
wire buttonA_debounced;
//Button B synchronisation and debouncing
wire buttonB_debounced;

//PSRAM interface
wire [15:0] data_out;      //Data read -> Output reg from PSRAM

//Reg
//PSRAM interface
//reg [23:0] address;      //Address of message to be written/read
reg [15:0] data_in;        //Data to be written (16 bits)
reg [15:0] read;           //Auxiliary Data read -> reg to be changed at procedural script
reg error;                 //Error flag

// Debugging
reg [3:0] proccess; //Keep track of write and reading test proccesses
reg [3:0] counter; //Counter to control debugging LEDs when pressing buttonA
reg pause;


//-----------------------------------------------------------------------------------------------------------------

//SUBMODULES

//84Mhz generated by Gowin's PLL
gowin_rpll_27_to_84 clk2(
    .clkout(clk_PSRAM), //84 MHz
    .clkin(sys_clk) //27MHz
);

//Debouncing proccesses to avoid noise from button pressing
sync_debouncer debuttonA(
    .clk(clk_PSRAM),
    .button(buttonA),
    .button_once(buttonA_debounced)
);
sync_debouncer debuttonB(
    .clk(clk_PSRAM),
    .button(buttonB),
    .button_once(buttonB_debounced)
);

//PSRAM initialization
psram initialize(
    //input
    .mem_clk(clk_PSRAM),
    .startbu(buttonB_debounced),
    .address(address),
    .read_write(read_write_uart),
    .data_in(data_in),

    //output
    .qpi_on(qpi_on),
    .endcommand(endcommand),
    .mem_ce(mem_ce),
    .data_out(data_out),
    .read_psram(read_psram),

    //inout
    .mem_sio(mem_sio),
    .message(message)
);

//UART1 channel communication
uart #(.DELAY_FRAMES(234), .BUFFER_LENGTH(BUFFER_LENGTH)) UART1 (
    //input
    .sys_clk(sys_clk),
    .uart_rx(uart_rx),
    .read_psram(read_psram),
    

    //output
    .read_write_uart(read_write_uart),
    .message(message),
    .address(address),
    .uart_tx(uart_tx)
);

//-----------------------------------------------------------------------------------------------------------------

//LOCAL PARAMETERS

//Testbench read & write
localparam [3:0] IDLE = 0;
localparam [3:0] DEBUG = 1;

//CHANGING PARAMETERS
localparam [15:0] ADDRESSA = 16'h01;
localparam [15:0] ADDRESSB = 16'h01;
localparam [15:0] MSGA = 16'h0121;
localparam [15:0] MSGB = 16'h0123;

//Number of bytes stored in buffer
localparam BUFFER_LENGTH = 6;

//-----------------------------------------------------------------------------------------------------------------

//SCRIPT

initial begin
    proccess <= 0;
    error <= 0;
    counter <= 0;
    pause <= 0;
end

always @(posedge clk_PSRAM) begin

   //DEBUGGING SECTION
   //Activates only when error is present while pressing buttonA
   if((error || proccess == DEBUG) && buttonA_debounced) begin

        counter <= counter + 1'd1;

        //For each button pressed, change debug leds

        case(counter) 
            0: led[3:0] <= read[15:12];
            1: led[3:0] <= read[11:8];
            2: led[3:0] <= read[7:4];
            3: led[3:0] <= read[3:0];
            4: begin
                led[3:0] <= 4'b1111;
                counter <= 0;

            end
            default: begin
                counter <= 0;
            end
        endcase
    end

    //Testing PSRAM communication
    if (qpi_on) begin  //if on IDLE state

      //White LED to begin proccess
      led_rgb[2:0] <= 3'b000;

      //LED RGBs
      if(error) led_rgb[2:0] <= 3'b011;           //Red LED
      else if (proccess == DEBUG) led_rgb[2:0] <= 3'b110;    //Blue LED = debugging state
      else led_rgb[2:0] <= 3'b101;    //Green LED = IDLE state, awaiting button
        
        case(pause)

          0: begin
            case (proccess)

              //Writing operation
              IDLE: begin
                if(endcommand && !read_psram) write <= message;
                if(endcommand && read_psram) begin
                    proccess <= DEBUG;
                    pause <= 1;
                end
              end

              //Awaits for instructions
               DEBUG: begin   
                 if (read == write) begin   
                    error <= 0; 
                  end
                  else error <= 1;
                  proccess <= IDLE;
               end
            endcase
          end
    
          1: begin //Awaits for button pressed
            if(buttonB_debounced) pause <= 0;
          end

        endcase
      end
end

endmodule

