//ReadMe: Top module for testing purposes.
//Refer to Testbench.v for simulation purposes
//PSRAM communication without the need to state beginning and ending of communication, but cant proccess same operations without a possible reset.
//-----------------------------------------------------------------------------------------------------------------

//Include sub-modules
//`include "PSRAM.v" //Simulation modules
//`include "gowin_rpll/grPLL_27_to_84.v" //rPLL Gowin native module

module TOP (

//IO pins
//INPUT
input sys_clk, //Internal 27 MHz oscillator
input buttonA, //Tang Nano Button A
input buttonB, //Tang Nano Button B

//PSRAM mem chip
inout wire [3:0] mem_sio,    // sio[0] pin 40, sio[1] pin 39, sio[2] pin 38, sio[3] pin 41
output mem_ce,               // pin 42
output clk_PSRAM,            // pin 6

//OUTPUT
//Debug RGB LED
output reg [2:0] led_rgb,             //RGB LEDs

//Debug external LEDs
output reg [3:0] led
);

//Variables
//Write/read variables
//Wire
wire [15:0] data_out;      //Data read -> wire cause it is output from PSRAM

//Reg
reg [23:0] address;        //Address of message to be written/read


wire [15:0] message;
reg [15:0] msg_reg = 0;


//assign message = (read_write == 0) ? msg_reg:16'hz;
assign message = (read_write == 1) ? msg_reg:16'hz;


reg [1:0] read_write;               //Read enable switch]
//reg read_write;               //Read enable switch
//  R   W   RW
//  0   0   0   :   Idle state
//  0   1   1   :   Writintg
//  1   0   2   :   Reading
//  1   1   3   :   Undefined
//reg quad_start;
reg [15:0] data_in;        //Data to be written (16 bits)
reg [15:0] read;           //Auxiliary Data read -> reg to be changed at procedural script
reg error;                 //Error flag

// Reg
reg [3:0] proccess; //Keep track of write and reading test proccesses
reg [3:0] counter; //Counter to control debugging LEDs when pressing buttonA
reg pause;

//Button A synchronisation and debouncing
wire buttonA_debounced;

//Button B synchronisation and debouncing
wire buttonB_debounced;


//84Mhz generated by Gowin's PLL
gowin_rpll_27_to_84 clk2(
    .clkout(clk_PSRAM), //84 MHz
    .clkin(sys_clk) //27MHz
);


//Debouncing proccesses to avoid noise from button pressing
sync_debouncer debuttonA(
    .clk(clk_PSRAM),
    .button(buttonA),
    .button_once(buttonA_debounced)
);

sync_debouncer debuttonB(
    .clk(clk_PSRAM),
    .button(buttonB),
    .button_once(buttonB_debounced)
);

//PSRAM initialization
psram initialize(
    //input
    .mem_clk(clk_PSRAM),
    .startbu(buttonB),
    .address(address),
    .read_write(read_write),
    //.quad_start(quad_start),
//    .data_in(data_in),


    //output
    .qpi_on(qpi_on),
    .endcommand(endcommand),
    .mem_ce(mem_ce),
//    .data_out(data_out),

    //inout
    .mem_sio(mem_sio),
    .message(message)
);

//Testbench read & write
localparam [3:0] WRITEA = 0;
localparam [3:0] WRITEB = 1;
localparam [3:0] READA = 2;
localparam [3:0] READB = 3;
localparam [3:0] WAITA = 4;
localparam [3:0] WAITB = 5;

//CHANGING PARAMETERS
localparam [15:0] ADDRESSA = 16'h01;
localparam [15:0] ADDRESSB = 16'h01;
localparam [15:0] MSGA = 16'h3547;
localparam [15:0] MSGB = 16'h9093;



initial begin
    proccess <= 0;
    error <= 0;
    //quad_start <= 0;
    counter <= 0;
    pause <= 0;
    read_write <= 0;
end

always @(posedge clk_PSRAM) begin

   //Activates only when error is present while pressing buttonA
   if((error || proccess == WAITA || proccess == WAITB) && buttonA_debounced) begin

        counter <= counter + 1'd1;

        //For each button pressed, change debug leds

        case(counter) 
            0: led[3:0] <= read[15:12];
            1: led[3:0] <= read[11:8];
            2: led[3:0] <= read[7:4];
            3: led[3:0] <= read[3:0];
            4: begin
                led[3:0] <= 4'b1111;
                counter <= 0;

            end
            default: begin
                counter <= 0;
            end
        endcase
    end

    //White LED to begin debugging
    led_rgb[2:0] <= 3'b000;

    //Testing PSRAM communication
    if (qpi_on) begin  //if on IDLE state

      //LED RGBs
      if(error) led_rgb[2:0] <= 3'b011;           //Red LED
      else if ((proccess == WAITA || proccess == WAITB)) led_rgb[2:0] <= 3'b110;    //Blue LED = waiting state
      else if ((proccess == WRITEA || proccess == WRITEB)) led_rgb[2:0] <= 3'b010;    //Blue LED = waiting state
      else if ((proccess == READA || proccess == READB)) led_rgb[2:0] <= 3'b001;    //Yellow LED = waiting state
      else led_rgb[2:0] <= 3'b111;    //LEDs off = Idle, awaiting button
        
        case(pause)

          0: begin
            case (proccess)

              //Writing operation
              WRITEA: begin   
                address <= ADDRESSA;
                msg_reg <= MSGA;
//                data_in <= MSGA;
                read_write <= 1;
                //read_write <= 0;
                //quad_start <= 1;
                if(endcommand) begin
                    proccess <= READA;
                    //quad_start <= 0;
                    //pause <= 1;
                end
              end

              //Reading operation
              READA: begin
                address <= ADDRESSA;
                read_write <= 2;
                //read_write <= 1;
                //quad_start <= 1;
                if(endcommand) begin 
                  proccess <= WAITA;
                  //quad_start <= 0;
                  //pause <= 1;
                  read <= message;
                  //read <= data_out;
                end
              end

              //Awaits for instructions
               WAITA: begin   
                 if ( read == MSGA ) begin   
                    error <= 0; 
                  end
                  else error <= 1;
                  proccess <= WRITEB;
               end

              //Writing operation
              WRITEB: begin   
                address <= ADDRESSB;
                msg_reg <= MSGB;
  //              data_in <= MSGB;
                read_write <= 1;
                //read_write <= 0;
                ////quad_start <= 1;
                if(endcommand) begin
                    proccess <= READB;
                    ////quad_start <= 0;
                    //pause <= 1;
                end
              end

              //Reading proccess
              READB: begin
                address <= ADDRESSB;
                read_write <= 2;
                //read_write <= 1;
                //quad_start <= 1;
                if(endcommand) begin 
                  proccess <= WAITB;
                  //quad_start <= 0;
                  //pause <= 1;
                  read <= message;
                  //read <= data_out;
                end
              end

              //Awaits for instructions
              WAITB: begin   
                 if ( read == MSGB ) begin   
                    error <= 0;
                    led_rgb[2:0] <= 3'b101;     //Comms' succeeded
                  end
                  else error <= 1;
               end
            endcase    
          end

          1: begin //Awaits for button pressed
            if(buttonB_debounced) pause <= 0;
          end

        endcase
      end
end

endmodule

