//ReadMe: Top module for testing purposes.
//Refer to Testbench.v for simulation purposes
//PSRAM communication WITH the need to state beginning and ending of communication. Choosen architecture due to future work (fingers crossed)
//-----------------------------------------------------------------------------------------------------------------

//Include sub-modules
//`include "PSRAM.v" //Simulation modules
//`include "gowin_rpll/grPLL_27_to_84.v" //rPLL Gowin native module

module TOP (

//IO pins
//INPUT
input sys_clk,                  //Internal 27 MHz oscillator
input buttonA,                  //Tang Nano Button A
input buttonB,                  //Tang Nano Button B

//PSRAM mem chip
inout [3:0] mem_sio,           // sio[0] pin 40, sio[1] pin 39, sio[2] pin 38, sio[3] pin 41
output mem_ce,                 // pin 42
output mem_clk_en,             // pin 6

//OUTPUT
//Debug RGB LED
output reg [2:0] led_rgb       //RGB LEDs

);

//Variables
//Write/read variables
wire [15:0] message;          // inout variable responsible to send and receive commands to be written and readen, respectively
wire quad_start;              // Flag to start QPI communication
wire [15:0] data_out;         // data output

//Reg
//PSRAM communication
reg [23:0] address;           // Address of message to be written/read
reg [15:0] msg_reg = 0;       // Reg variable of message used in procedural assignment
reg com_start;                // Register - indicates whether start QPI or not
reg d_com_start;              // Register - stores com_start value to detect step-up

reg [1:0] read_write;         // Read enable switch
//  R   W   RW
//  0   0   0   :   Idle state
//  0   1   1   :   Writintg
//  1   0   2   :   Reading
//  1   1   3   :   Undefined

//DEBUGGING
reg [15:0] read;            //Auxiliary Data read -> reg to be changed at procedural script -> debug LEDs
reg error;                  //Error flag
reg [3:0] counter;          //Counter to control debugging LEDs when pressing buttonA
reg pause;                  //Pause flag in order to debug. Proccess MUST work without pauses

//TOP operation
reg [3:0] proccess;         //Keep track of write and reading test proccesses
reg [15:0] data_in;

//Rising edge
assign quad_start = (com_start & ~d_com_start);

//Button A synchronisation and debouncing
wire buttonA_debounced;

//Button B synchronisation and debouncing
wire buttonB_debounced;

//84Mhz generated by Gowin's PLL
gowin_rpll_27_to_84 clk2(
    .clkout(clk_PSRAM), //84 MHz
    .clkin(sys_clk) //27MHz
);

//Debouncing proccesses to avoid noise from button pressing
sync_debouncer debuttonA(
    .clk(clk_PSRAM),
    .button(buttonA),
    .button_once(buttonA_debounced)
);

sync_debouncer debuttonB(
    .clk(clk_PSRAM),
    .button(buttonB),
    .button_once(buttonB_debounced)
);

//PSRAM initialization
psram initialize(
    //input
    .mem_clk(clk_PSRAM),
    .startbu(buttonB),
    .address(address),
    .read_write(read_write),
    .quad_start(quad_start),
    .data_in(data_in),

    //output
    .mem_clk_en(mem_clk_en),
    .qpi_on(qpi_on),
    .endcommand(endcommand),
    .mem_ce(mem_ce),
    .data_out(data_out),

    //inout
    .mem_sio(mem_sio),
    .message(message)
);

//Testbench read & write
localparam [3:0] WRITEA = 0;
localparam [3:0] WRITEB = 1;
localparam [3:0] READA = 2;
localparam [3:0] READB = 3;
localparam [3:0] WAITA = 4;
localparam [3:0] WAITB = 5;

//CHANGING PARAMETERS
//localparam [22:0] ADDRESSA = 23'h7FFFFF;
localparam [22:0] ADDRESSA = 23'h7FFFFE;
localparam [15:0] ADDRESSB = 16'hABCD;
localparam [15:0] MSGA = 16'h1234;
localparam [15:0] MSGB = 16'h4464;

// Declaração de variáveis auxiliares
integer i;                  // Loop iteration
integer erro_data_out;      // Data_out error
integer erro_read;          // Read error
reg [15:0] rand_data;       // Random data_in

// Pseudorandom 16-bits LFSR
reg [15:0] lfsr;

// Pseudorandom 4-bits LFSR
reg [3:0] lfsr_a;  // Primeira parte do LFSR
reg [3:0] lfsr_b;  // Segunda parte do LFSR
reg [3:0] lfsr_c;  // Terceira parte do LFSR
reg [3:0] lfsr_d;  // Quarta parte do LFSR

initial begin
    proccess <= WRITEA;
    error <= 0;
    counter <= 0;
    pause <= 0;
    read_write <= 0;
    com_start <= 0;
    d_com_start <= 0;
    read <= 16'hffff;
    address <= 22'h0000;
    i <= 0;
    rand_data <= 0;
    erro_data_out <= 0;
    erro_read <= 0;
    lfsr <= 16'hAFAF;  // Seed inicial para o LFSR
    led_rgb <= 4'b0000;
    lfsr_a <= 4'hf;  // Seed inicial para o LFSR A
    lfsr_b <= 4'hf;  // Seed inicial para o LFSR B
    lfsr_c <= 4'hf;  // Seed inicial para o LFSR C
    lfsr_d <= 4'hf;  // Seed inicial para o LFSR D
end

always @(posedge clk_PSRAM) begin

    led_rgb <= 4'b110;

    d_com_start <= com_start;

    lfsr <= {lfsr[14:0], lfsr[15] ^ lfsr[13] ^ lfsr[12] ^ lfsr[10]};
    // Atualiza cada LFSR individualmente, com taps diferentes para cada um
    lfsr_a = {lfsr_a[2:0], lfsr_a[3] ^ lfsr_a[2]};  // LFSR A (tap positions 3 e 2)
    lfsr_b = {lfsr_b[2:0], lfsr_b[3] ^ lfsr_b[1]};  // LFSR B (tap positions 3 e 1)
    lfsr_c = {lfsr_c[2:0], lfsr_c[3] ^ lfsr_c[2] ^ lfsr_c[1]};  // LFSR C (tap positions 3, 2 e 1)
    lfsr_d = {lfsr_d[2:0], lfsr_d[3] ^ lfsr_d[0]};  // LFSR D (tap positions 3 e 0)

    if (qpi_on) begin

            led_rgb <= 4'b000;
        case (proccess)
            WRITEA: begin
                // Incrementa o endereço e gera dados aleatórios
                if (i <= 23'h7FFFFF) begin
                    //if(!com_start) rand_data = lfsr; //Se a comunicação não tiver começado, atribui um valor pseudo-aleatório para rand_data, que será utilizado como critério de erros.
                    if (!com_start) begin
                        //rand_data = 16'hFEFE;
                        // Combina os 4 LFSRs em um valor final de 16 bits
                        rand_data = {lfsr_a, lfsr_b, lfsr_c, lfsr_d};  // Concatena os LFSRs
                        //rand_data = lfsr[15:0];
                        data_in = rand_data;  // Gera dados aleatórios de 16 bits
                    end
                    address <= i[22:0];  // Atribui o valor do endereço
                    read_write <= 1;  // Sinaliza operação de escrita
                    com_start <= 1;

                    if (endcommand) begin
                        proccess <= READA;
                        com_start <= 0;
                    end
                end
            end

            READA: begin
                // Lê os dados no mesmo endereço
                read_write <= 2;  // Sinaliza operação de leitura
                com_start <= 1;

                if (endcommand) begin
                    read <= data_out;  // Armazena o valor lido
                    com_start <= 0;
                    proccess <= WAITA;
                end
            end

            WAITA: begin
                // Compara o valor lido com o valor escrito
                if (read != rand_data) begin
                    error <= 1;  // Acusa erro se os valores forem diferentes
                    erro_read <= erro_read + 1;
                    //data_aux <= read;  // Armazena o valor lido incorreto
                end
                if (data_out != rand_data) begin
                    error <= 1;
                    erro_data_out <= erro_data_out + 1;
                end

                if (error) begin
                    error <= 1;  // Reseta a flag de erro
                end

                // Incrementa o endereço em 2, pois cada escrita/leitura compreende 2 bytes de memória
                i = i + 2;

                // Se atingir o limite de endereço, termina
                if (i >= 23'h7FFFFF) begin
                    proccess <= WAITB;
                end
                else begin
                    proccess <= WRITEA;  // Continua o processo de escrita/leitura
                end
            end

            WAITB: begin
                proccess <= WAITB;
                // Verificação final de status
                if (!error) begin
                    led_rgb[2:0] <= 3'b101;  // Sucesso
                end
                else begin
                    led_rgb[2:0] <= 3'b011;  // Indica erro
                end
            end
        endcase
    end
end
endmodule

