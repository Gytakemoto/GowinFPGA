//ReadMe: Top module for testing purposes.
//Refer to Testbench.v for simulation purposes
//-----------------------------------------------------------------------------------------------------------------

//Include sub-modules
//`include "PSRAM.v" //Simulation modules
//`include "gowin_rpll/grPLL_27_to_84.v" //rPLL Gowin native module

module TOP (

//IO pins
//INPUT
input sys_clk, //Internal 27 MHz oscillator
input buttonA, //Tang Nano Button A
input buttonB, //Tang Nano Button B

//PSRAM mem chip
inout wire [3:0] mem_sio,    // sio[0] pin 40, sio[1] pin 39, sio[2] pin 38, sio[3] pin 41
output mem_ce,               // pin 42
output clk_PSRAM,            // pin 47

//OUTPUT
//Debug RGB LED
output reg [2:0] led_rgb,             //RGB LEDs
//led_rgb[2]: RED LED pin 9
//led_rgb[1]: GREEN_LED pin 11
//led_rgb[0]: BLUE_LED pin 10

//Debug external LEDs
output reg [3:0] led
);

//Variables

//Write/read variables
//Wire
wire [15:0] data_out;      //Data read -> wire cause it is output from PSRAM

//Reg
reg [23:0] address;        //Address of message to be written/read
reg write_sw;              //Write enable switch
reg read_sw;               //Read enable switch
reg [15:0] data_in;        //Data to be written
reg [15:0] read;           //Auxiliary Data read -> reg to be changed at procedural script
reg error;                 //Error flag

// Reg
reg [3:0] estepe; //APAGAR depois
reg [3:0] counter; //Counter to control debugging LEDs when pressing buttonA
reg pause;

//Button A synchronisation and debouncing
wire buttonA_synched;
wire buttonA_debounced;

//84Mhz generated by Gowin's PLL
gowin_rpll_27_to_84 clk2(
    .clkout(clk_PSRAM), //84 MHz
    .clkin(sys_clk) //27MHz
);

//Button A sync and debouncer
sync sync_buttonA(
    .clock(clk_PSRAM),
    .in(buttonA),
    .out(buttonA_synched)
);

debouncer deb_buttonA(
    .clock(clk_PSRAM),
    .in(buttonA),
    .out(buttonA_debounced)
);

//PSRAM initialization
psram initialize(
    //input
    .mem_clk(clk_PSRAM),
    .startbu(buttonB),
    .address(address),
    .read_sw(read_sw),
    .write_sw(write_sw),
    .data_in(data_in),

    //output
    .qpi_on(qpi_on),
    .endcommand(endcommand),
    .mem_ce(mem_ce),
    .data_out(data_out),

    //inout
    .mem_sio(mem_sio)
);

//Testbench read & write
localparam [3:0] WRITEA = 0;
localparam [3:0] WRITEB = 1;
localparam [3:0] READA = 2;
localparam [3:0] READB = 3;
localparam [3:0] NEXT = 4;

initial begin
    estepe <= 0;
    error <= 0;
    write_sw <= 0;
    read_sw <= 0;
    counter <= 0;
end

function button_pressed(button);

  reg [15:0] sync_button;

  begin
  sync_button = {sync_button[2:0],button};
  button_pressed = ~sync_button[3] & sync_button[2];
  end  
endfunction

always @(posedge clk_PSRAM) begin

   //Activates only when error is present while pressing buttonA
   if(error && !buttonA_debounced) begin

        counter <= counter + 1'd1;

        //For each button pressed, change debug leds

/*
        case(counter) 
            0: led[3:0] <= data_out[15:12];
            1: led[3:0] <= data_out[11:8];
            2: led[3:0] <= data_out[7:4];
            3: led[3:0] <= data_out[3:0];
            //4: led[3:0] <= 4'b1001;
            default: begin
                counter <= 0;
            end
        endcase
*/
/*
         case(counter) 
            0: led[3:0] <= 4'b0000;
            1: led[3:0] <= 4'b0010;
            2: led[3:0] <= 4'b0011;
            3: led[3:0] <= 4'b0100;
            4: led[3:0] <= 4'b0101;
            default: begin
                counter <= 0;
            end
        endcase
*/

        led[3:0] <= counter;
        
        if(counter >= 4'd15) counter <= 0;
    end

  //LED RGBs
  if(error) led_rgb[2:0] <= 3'b011;           //Red LED
  else if (!pause) led_rgb[2:0] <= 3'b110;     //Blue LED = Proccessing
  else if (qpi_on && pause) led_rgb[2:0] <= 3'b101;    //Green LED = Idle, awaiting button


    //Testing PSRAM communication
    if (qpi_on && !error) begin  //if on IDLE state
        
        case(pause)

          0: begin
            case (estepe)
              WRITEA: begin   
                address <= 8'hFA;
                data_in <= 16'h1234;
                write_sw <= 1;
                if(endcommand) begin
                    estepe <= WRITEB;
                    write_sw <= 0;
                    pause <= 1;
                end
              end
              WRITEB: begin   
                address <= 8'h2;
                data_in <= 16'h5678;
                write_sw <= 1;
                if(endcommand) begin
                    estepe <= READA;
                    write_sw <= 0;
                    pause <= 1;
                end
              end
              READA: begin
                address <= 8'hFA;
                read_sw <= 1;
                if(endcommand) begin 
                  estepe <= READB;
                  read_sw <= 0;
                  pause <= 1;
                end
              end
              READB: begin
                read <= data_out;
                if ( data_out != 16'h1234 ) begin   
                  error <= 1; 
                end
                address <= 8'h2;
                read_sw <= 1;
                if(endcommand) begin 
                  estepe <= NEXT;
                  read_sw <= 0;
                  pause <= 1;
                end
              end
              /*
              NEXT: begin
                read <= data_out;
                if ( data_out != 16'h5678 ) begin 
                  error <= 1;
                end
                //if(endcommand) estepe <= WRITEA;
              end   
*/     
            endcase    
          end

          1: begin //Awaits for button pressed
            if(!buttonB) pause <= 0;
          end

        endcase
      end
end

endmodule

