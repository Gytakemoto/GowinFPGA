
/* ------------------------------- TOP MODULE ------------------------------- */
module TOP (

//Tang Nano 1k
input sys_clk,                	// Internal 27 MHz oscillator

//UART
input uart_rx,                 	// RX UART wire [pin 18]

//Data acquisition
input buttonA, 					//Button that requests data acquisition		

//PSRAM mem chip
inout [3:0] mem_sio,     		// Communication busbar for PSRAM communication - [sio[0] pin 40, sio[1] pin 39, sio[2] pin 38, sio[3] pin 41]
output mem_ce,                	// PSRAM chip enable - [pin 42]
output mem_clk_enabled,         // PSRAM clock pin - [pin 6]
output uart_tx,                	// TX UART wire [pin 17]

//DEBUGGING
//Debug RGB LED
output reg [2:0] led_rgb     	// RGB LEDs
);

/* -------------------------------- Variables ------------------------------- */

/* ----------------------------- PSRAM interface ---------------------------- */

// Inputs (from PSRAM.v module)
wire clk_PSRAM;				   // 84MHz rPLL generated clock. Used in PSRAM interface
//wire endcommand;			   // Input flag - indicates whether PSRAM writing or reading finished
wire qpi_on;				   // Input flag - indicates whether QPI communication is on

// Outputs (to PSRAM.v module) - Determined by "MCU" or UART
//reg [22:0] address;       	   // Address of message to be written/read
//reg [15:0] data_in;            // Data to be written (16 bits)
reg [15:0] read;               // Auxiliary Data read -> reg receives data_out in a procedural script
wire [15:0] data_out;      	   // Data read -> Output reg from PSRAM
//reg [1:0] read_write;		   // Define read or write proccess
	//read_write
	//0	0 : Do nothing
	//0	1 : Write data from PSRAM
    //1	0 : Read data to PSRAM
    //1	1 : Do nothing


/* ----------------------------- UART interface ----------------------------- */

// Inputs (from UART.v module)
	// Request read or write through UART
//wire quad_start_uart;         // Start reading OR writing proccess via UART
//wire [1:0] read_write_uart;   // Read or write switch via UART
//wire [22:0] address_uart;     // Address of interest (write or read) via UART
//wire [15:0] data_in_uart;     // Data to be written via UART

wire [7:0] threshold;             // Threshold type: "T" or "B"]
wire [23:0] samples_after;        // Number of samples to be written after the threshold
wire [23:0] samples_before;       // Number of samples to be written before the threshold
wire start_acq;				//Flag to start acquisition
reg [1:0] read_write_acq;
reg [22:0] address_acq;
reg [15:0] data_in_acq;

// Outputs (to UART.v module)
reg send_uart;				  // Flag - inform UART to send data through Tx

/* -------------------------- Internal variables -------------------------- */

reg error;                  // Error flag
reg [3:0] process; 			// State-machine of top.v states

// Request read or write through MCU
reg com_start;				// Detect rising edge to start quad_start
reg d_com_start;			
reg quad_start;            	// Output flag - Start reading OR writing proccess via MCU
	// quad_start = com_start && !d_com_start;

// Directly control write and read process, through MCU (Gowin)
reg quad_start_mcu;
reg [1:0] read_write_mcu;
reg [22:0] address_mcu;
reg [15:0] data_in_mcu;
reg [1:0] read_write;
reg [22:0] address;
reg [15:0] data_in;



/* ----------------------- Data acquisition interface ----------------------- */

reg [22:0] i;
reg [22:0] i_pivot; 			//Refers to the sample where threshold was detected
reg [22:0] i_pivot_valid;
reg [22:0] address_debug;
reg [22:0] new_address;	
reg d_flag_acq;
wire flag_acq;
reg start_acquisition;
reg [1:0] buttons_pressed;			//Number of times the buttonA was pressed
reg [11:0] adc_data_in;				//Simulates 12-bit adc data
reg stop_acquisition;
reg condition1;
reg condition2;
reg condition3;
reg condition_met;

wire [22:0] i_minus_i_pivot = i - i_pivot;
wire [22:0] i_max_minus_i_pivot_plus_i = i_max - i_pivot + i;
reg [22:0] i_minus_i_pivot_reg;
reg [22:0] samples_after_adjusted;
reg condition1_reg, condition2_reg, condition3_reg;

/* ------------------------------- Submodules ------------------------------- */

/* --------------------- 84Mhz generated by Gowin's PLL --------------------- */
gowin_rpll_27_to_84 clk2(
	.clkout(clk_PSRAM), 	// 84 MHz
	.clkin(sys_clk) 		// 27MHz
);

/* ---------------------------------- PSRAM --------------------------------- */
psram initialize(
	//input
	.mem_clk(clk_PSRAM),
	.address(address_mcu),
	.read_write(read_write_mcu),
	.data_in(data_in_mcu),
	.quad_start(quad_start_mcu),

	//output
	.mem_clk_enabled(mem_clk_enabled),
	.qpi_on(qpi_on),
	.endcommand(endcommand),
	.mem_ce(mem_ce),
	.data_out(data_out),

	//inout
	.mem_sio(mem_sio)
);

/* ----------------------- UART1 channel communication ---------------------- */
uart #(.DELAY_FRAMES(729), .BUFFER_LENGTH(BUFFER_LENGTH)) UART1 (
	//input
	.clk_PSRAM(clk_PSRAM),
	.uart_rx(uart_rx),
	.send_msg(read),
	.send_uart(send_uart),
	
	//output
	//.led(led),
	//.read_write(read_write_uart),
	//.quad_start(quad_start_uart),
	//.data_in(data_in_uart),
	//.address(address_uart),

	.threshold(threshold),
    .samples_after(samples_after),        // Number of samples to be written after the threshold
    .samples_before(samples_before),       // Number of samples to be written before the threshold
    .flag_acq(flag_acq), 

	.uart_tx(uart_tx)
);

/* ---------------------------- Local parameters ---------------------------- */

//Testbench read & write
localparam [3:0] WRITE_MCU_INIT = 0;
localparam [3:0] READ_MCU_INIT = 1;
localparam [3:0] CHECK_STARTUP = 2;
localparam [3:0] IDLE = 3;
localparam [3:0] DATA_ACQUISITION = 4;

//Maximum number of 2-byte addresses (12-bit samples): 8 MB / 2 = 4 MB
//Same as 2^22 = 4MB
//PSARM has 23 bits for addressing, which means that it supports the maximum address # of 8.388.608 - 1 = 8.388.607
//The maximum iteration must be at 2^22 = 4.194.304:
//() * 2 = 8.388.606; thus in the last iteration it will write in the 8.388.606 and 8.388.607
localparam [22:0] i_max = 1 << 22;

//Buffer's bytes length
localparam BUFFER_LENGTH = 10;

/* ---------------------------- Button debouncing --------------------------- */

//Button A synchronisation and debouncing
wire buttonA_debounced;

//Debouncing proccesses to avoid noise from button pressing

sync_debouncer debuttonA(
    .clk(clk_PSRAM),
    .button(buttonA),
    .button_once(buttonA_debounced)
);

/* --------------------------- Procedural routine --------------------------- */

initial begin
	process <= WRITE_MCU_INIT;
	error <= 0;
	read <= 0;
	send_uart <= 0;
	com_start <= 0;
	d_com_start <= 0;

	//MCU read-write variables
	read_write_mcu <= 0;
	address_mcu <= 22'hzzzz;
	data_in_mcu <= 0;
	quad_start_mcu <= 0;
    led_rgb <= 3'b111;

	//Acquisition variables
	i_pivot = 0;
    start_acquisition = 0;
    buttons_pressed <= 0;
	stop_acquisition <= 0;
	address_debug <= 0;
end

always @(posedge clk_PSRAM) begin     
	//* Constantly update regulators in order to avoid inferred latches
	/*
    quad_start <= 0;
	read_write <= read_write;
	address <= address;
	data_in <= data_in;
	read <= read;
	send_uart <= 0;
    */
	// Detect a rising edge of mcu requisition. Only valid on MCU controlling of WRITE/READs
	quad_start_mcu <= (com_start && ~d_com_start);
	d_com_start <= com_start;
	com_start <= 0;

	// Detect a rising edge of UART requisition
	start_acquisition <= (flag_acq && ~d_flag_acq);
	d_flag_acq <= flag_acq;


    // Routine to detect source of requisition: UART or MCU
	if(quad_start_mcu) begin
        if(process == DATA_ACQUISITION) begin
            read_write <= read_write_acq;
            address <= address_acq;
            data_in <= data_in_acq;
            quad_start <= quad_start_mcu;
        end
        else begin
        read_write <= read_write_mcu;
        address <= address_mcu;
        data_in <= data_in_mcu;
        quad_start <= quad_start_mcu;
        end
    end



// if else if else is bad

	//* Only when QPI is ready
	if (qpi_on) begin
		case (process)
		//todo: inserir uma verificação de aquisição fora do IDLE
		//todo: semelhante ao todo lá embaixo, talvez expandido para qualquer fluxo na implementação final
		    // Writing operation to test PSRAM before starting
			WRITE_MCU_INIT: begin
				address_mcu <= 24'hABCD;
				data_in_mcu <= 16'h1234;
				read_write_mcu <= 1;
				com_start <= 1;
				if(endcommand) begin
					com_start <= 0;
					process <= READ_MCU_INIT;
				end
			end
			READ_MCU_INIT: begin
				address_mcu <= 24'hABCD;
				read_write_mcu <= 2;
				com_start <= 1;
				if(endcommand) begin
					read <= data_out;
					read_write_mcu <= 0;
					com_start <= 0;
					process <= CHECK_STARTUP;
				end
			end
			CHECK_STARTUP: begin
				//* If writing and reading processess were OK
				if(read == data_in_mcu) begin
					led_rgb <= 3'b101;
					error <= 0;
					process <= IDLE;
				end
				// If not...
				else begin
                    led_rgb[2:0] <= 3'b011;
					error <= 1;
				end
			end

			IDLE: begin
				
				//Start acquisition rising edge detected
				if(start_acquisition) begin
					process <= DATA_ACQUISITION;
					//* Always begin from start
					i <= 1;						//First sample -> 0 address
					buttons_pressed <= 0;		//Reset threshold button
					i_pivot = 0;				//Reset pivot
					adc_data_in <= 0;
					stop_acquisition <= 0;
                    led_rgb[2:0] <= {led_rgb[2:0] + 3'd1};
				end else process <= IDLE;

			end
			DATA_ACQUISITION: begin
			//todo: inserir um erro caso o processo ainda não esteja finalizado e outra aquisição seja requisitada pela ESP32
			//todo: pensei em:
			//todo: if(start_acquisition) led <= 3'b010; //Purple light if a data recquisition occurs during DATA_ACQUISITION process

				
				//*Validar button_debounced
                
				if(!buttonA_debounced) begin
					buttons_pressed <= buttons_pressed + 1'd1;
                    //When pressing for the first time, "detect threshold"
                    //todo: Incluir uma condição para verificar se o tipo de requisição é por botão
                end
                if(buttons_pressed == 1'd1) begin
                        i_pivot = i;
                        i_pivot_valid = 1;
                        address_debug <= i_pivot[22:0];
				end


				if(i < i_max) begin
					//If i_pivot = 0, it means threshold wasn't reached

                    //Caminho critico!!!!!!!

                    if (i_pivot_valid) begin
                        // Precompute intermediate values
                        i_minus_i_pivot_reg <= i - i_pivot;
                        samples_after_adjusted <= samples_after - (i_max - i_pivot);

                        // First stage: compute conditions
                        condition1_reg <= (samples_after == 23'd0);
                        condition2_reg <= (i >= i_pivot) && (i_minus_i_pivot_reg >= samples_after);
                        condition3_reg <= (i >= samples_after_adjusted);

                        // Second stage: compute final result
                        stop_acquisition <= (condition1_reg || condition2_reg || condition3_reg);
                    end

                    //todo: changed delay due to pipeline. Need to verify if logic's changed

					//While stop wasn't requested, write in memory
					if(!stop_acquisition) begin
							//12 bits fit in 16 bits						
							data_in_acq <= {4'b0000,adc_data_in};
							//address increases by 2 each time the sample updates
							//address starts from 0
							//!Same as: address_mcu <= 23'd2 *(i[21:0]-23'd1);

                            //todo: o acréscimo de um new_address causou um delay de um clock para a atribuição do address... CONSERTAR
                            new_address <= (i[22:0] - 23'd1) << 1;
							address_acq <= new_address;
							//@i_max:
							// address_mcu <= (2^22-1) * 2 = 8.388.606
							// then, it'll write 8.388.606 and 8.388.607
							read_write_acq <= 1;	//write in memory
							com_start <= 1;
							if(endcommand) begin
								com_start <= 0;
								//+1 for each iteration
								adc_data_in <= adc_data_in + 1'd1;
								i <= i + 1;		
							end
					end
					else begin
						read <= 16'hABCD;	//Dummy mesage to be read by ESP32
                        //led_rgb[2:0] <= {led_rgb[2:0] + 3'd1};
						send_uart <= 1;  	// Flag to send message via UART
						process   <= IDLE;   // After finishing the acquisition, go back to IDLEfter finishing the acquisition, go back to IDLE
					end
				end else i <= 1;			//Resetting number of samples to loop through PSRAM




			end

		endcase
	end
end
endmodule

